//  **************************************************
//  *              notif1 table design               *
//  **************************************************


module notif1_gate(input a, output y);
  assign y = ~a;
endmodule